import TestBenchTemplates::*;
import ministFifo::*;

//////////////////////////
// Functional Testbenches

// These testbenches compare the outputs of the fifo against a reference fifo.
// If there is any mismatch in the outputs, the simulator will print out an
// error message.

(* synthesize *)
module mkTbPipelineFunctional();
    Fifo#(Bit#(8)) fifo <- mkMyPipelineFifo();
    let m <- mkTbFunctionalTemplate(fifo, Pipeline);
endmodule


(* synthesize *)
module mkTbBypassFunctional();
    Fifo#(Bit#(8)) fifo <- mkMyBypassFifo();
    let m <- mkTbFunctionalTemplate(fifo, Bypass);
endmodule

(* synthesize *)
module mkTbCFFunctional();
    Fifo#(Bit#(8)) fifo <- mkMyCFFifo();
    let m <- mkTbFunctionalTemplate(fifo, CF);
endmodule


//////////////////////////
// Scheduling Testbenches

// These testbenches force the scheduling constraints that should be valid for
// each FIFO. These constraints include:
//
//  if the FIFO has an implemented clear method:
//      Bypass, CF:   {notFull, enq} < {notEmpty, first, deq} < clear
//      Pipeline, CF: {notEmpty, first, deq} < {notFull, enq} < clear
//  if the FIFO doesn't have an implemented clear method:
//      Bypass, CF:   {notFull, enq} < {notEmpty, first, deq}
//      Pipeline, CF: {notEmpty, first, deq} < {notFull, enq}
//
// If you get a compiler error while compiling any of these testbenches, then
// the FIFO does not meet the required scheduling constraints.

// Why don't you have to instantiate mkMyCFFifo before passing it to
// mkTbSchedulingTemplate? This testbench template takes a module constructor,
// not an interface. This testbench uses the module constructor to construct
// two copies of the same fifo for scheduling tests.

(* synthesize *)
module mkTbPipelineScheduling();
    let m <- mkTbSchedulingTemplate(mkMyPipelineFifo, Pipeline);
endmodule


(* synthesize *)
module mkTbBypassScheduling();
    let m <- mkTbSchedulingTemplate(mkMyBypassFifo, Bypass);
endmodule

(* synthesize *)
module mkTbCFScheduling();
    let m <- mkTbSchedulingTemplate(mkMyCFFifo, CF);
endmodule

